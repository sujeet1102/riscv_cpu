/*
# Author:		Sujeet Jagtap
# Module:		alu
# Description:	
# Inputs:		
# Outputs:		
*/
module alu (
	
);



endmodule